Architecture behavior of ej_combinacional_testbench is

   Component Ejercicio1 
	   Port(
		 SW1 : in STD_LOGIC;
		 SW2 : in STD_LOGIC;
		 LED : out STD_LOGIC);
	End component;
	
	
	signal SW1 : std_logic :='0';
	signal SW2 : std_logic :='0';

	signal LED : std_logic;
	
Begin 
   uut: Ejercicio1 port map (
	   SW1 => SW1,
		SW2 => SW2,
		LED => LED
	);
	
	stim_proc : process 
	begin 
	   SW1 <= '0'; SW2 <= '0'; wait for 10ns;
		SW1 <= '0'; SW2 <= '1'; wait for 10ns;
		SW1 <= '1'; SW2 <= '0'; wait for 10ns;
		SW1 <= '1'; SW2 <= '1'; wait for 10ns;
	wait;
	end process;
	end;