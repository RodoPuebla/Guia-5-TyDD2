library verilog;
use verilog.vl_types.all;
entity Ejercicio1_vlg_vec_tst is
end Ejercicio1_vlg_vec_tst;
