library verilog;
use verilog.vl_types.all;
entity Ejercicio1_vlg_check_tst is
    port(
        LED             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Ejercicio1_vlg_check_tst;
